module Strings;
 string s1="good";
  string s2="bad";
  string s3="ugly";
  string s4,s5,s6;
  initial begin
  s4="better";
  s5="worse";
    s6="";
    
    $display("s1=%s,s2=%s,s3=%s,s4=%s,s5=%s,s6=%s",s1,s2,s3,s4,s5,s6);
  end
endmodule

